
// alu function bits
//`define Fsize  1

`define RADD  1'b0
`define RMUL 1'b1
